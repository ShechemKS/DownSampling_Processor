module top_processor(	input wire clock, 				
								input wire start_process,
								output wire s0, s1, s2, s3,
								output endProcess);
								
								
								
	// For processor 
	wire [19:0] cm_out;						
	wire [7:0] dm_processor;				
	wire [31:0] im_out;						
	wire [1:0] status;						
	wire dm_r, dm_wr, cm_r, im_r;			
	wire [7:0] ac_out;						
	wire [9:0] pc_out;
	
	wire [2:0] mar_cm;						
	wire [19:0] mar_dm;						
	wire end_process;
	wire slow_clk;
		
	assign endProcess = end_process;	
					 
	// Main Controller

	
	// Memory DRAM
	
	wire [7:0] data_in_com; 				// data to the com module to be transmitted 
	wire [7:0] dm_in;							// data to the dram
	wire [7:0] dm_out;
	
	// Muxes
	wire [19:0] tx_dm;						// address from transmitter module to write
	wire [19:0] dm_addr;						// data memory address ( from processor or from tx_addr)
	wire [19:0] rx_dm;
	
	// Tx and Rx
	wire [7:0] dm_transmitter; 
	wire tx_en; 
	wire tx_clk_en, rx_clk_en;
	
	//wire tx, tx_busy; 
	wire [7:0] tx_data;
	wire [7:0] data_out_rx;					// data from receiver module
	
	

	C_ram 		cram1(.address(mar_cm),
							.clock(clock),
							.rden(cm_r),
							.q(cm_out));	
							
	iram  		iram1(	.clock(clock), 
								.im_r(im_r), 
								.addr(pc_out), 
								.instr_out(im_out)); 
					
	Processor 	cpu (		.clock(clock), 
								.cm_out(cm_out), 
								.dm_out(dm_processor), 
								.im_out(im_out), 
								.status(status), 
								.dm_r(dm_r), 
								.im_r(im_r), 
								.cm_r(cm_r), 
								.dm_wr(dm_wr), 
								.dm_in(ac_out), 
								.pc_out(pc_out), 
								.mar_dm(mar_dm), 
								.mar_cm(mar_cm),
								.end_process(end_process));
								
	dram	d_ram( 	.address(mar_dm),
						.clock(clock),
						.data(ac_out),
						.wren(dm_wr),
						.rden(dm_r), 
						.q(dm_processor));					

	main_control mc1(		.clock(clock), 
								.start_process(start_process),
								.end_process(end_process), 
								.status(status), 
								.s0(s0), .s1(s1), .s2(s2), .s3(s3)); 
			
	slowclock clk1 (	.inclk(clock),
							.outclk(slow_clk),
							.switch_clock(status));

					
endmodule 	
	
