module iram(	input clock, im_r,
					input [9:0] addr,
					output wire [31:0] instr_out);
	
	reg [31:0] memory [128:0];
	reg [31:0] current_instruction;
	
	initial begin
		//$readmemb("Inst_mem.mem", memory);
    memory[0]   = 32'b00100111110000000000000000000000;
    memory[1]   = 32'b00111000000000000000000000000011;
    memory[2]   = 32'b01100100100000000000000000000000;
    memory[3]   = 32'b00111000000000000000000000000100;
    memory[4]   = 32'b01100101000000000000000000000000;
    memory[5]   = 32'b00111000000000000000000000000101;
    memory[6]   = 32'b01100010100000000000000000000000;
    memory[7]   = 32'b00111000000000000000000000000110;
    memory[8]   = 32'b11110101100000000000000000000010;
    memory[9]   = 32'b01100011000000000000000000000000;
    memory[10]   = 32'b01010000000000000000000000000000;
    memory[11]   = 32'b00110000000000000000000000000000;
    memory[12]   = 32'b01100010000000000000000000000000;
    memory[13]   = 32'b10000000100000000000000000000000;
    memory[14]   = 32'b00110000000000000000000000000000;
    memory[15]   = 32'b10110000000000000000000000000000;
    memory[16]   = 32'b10011101101000000000000000000000;
    memory[17]   = 32'b01100010000000000000000000000000;
    memory[18]   = 32'b10000000100000000000000000000000;
    memory[19]   = 32'b00110000000000000000000000000000;
    memory[20]   = 32'b10011101101000000000000000000000;
    memory[21]   = 32'b10100000000000000000000000000000;
    memory[22]   = 32'b10100000000000000000000000000000;
    memory[23]   = 32'b11000110001010100000000000100001;
    memory[24]   = 32'b01011000000000000000000000000000;
    memory[25]   = 32'b01000000000000000000000000000000;
    memory[26]   = 32'b10000111000000000000000000000000;
    memory[27]   = 32'b11000111001100100000000000011101;
    memory[28]   = 32'b11000000000000000000000000001010;
    memory[29]   = 32'b10000001000000000000000000000000;
    memory[30]   = 32'b10000001000000000000000000000000;
    memory[31]   = 32'b00100100000000000000000000000000;
    memory[32]   = 32'b11000000000000000000000000001010;
    memory[33]   = 32'b01011000000000000000000000000000;
    memory[34]   = 32'b01000000000000000000000000000000;
    memory[35]   = 32'b01110101000000000000000000000000;
    memory[36]   = 32'b01100010100000000000000000000000;
    memory[37]   = 32'b00111000000000000000000000000100;
    memory[38]   = 32'b01100100100000000000000000000000;
    memory[39]   = 32'b00111000000000000000000000000011;
    memory[40]   = 32'b01100101000000000000000000000000;
    memory[41]   = 32'b11000000000000000000000000101010;
    memory[42]   = 32'b01010000000000000000000000000000;
    memory[43]   = 32'b00110000000000000000000000000000;
    memory[44]   = 32'b01100010000000000000000000000000;
    memory[45]   = 32'b10011110001100000000000000000000;
    memory[46]   = 32'b00110000000000000000000000000000;
    memory[47]   = 32'b10110000000000000000000000000000;
    memory[48]   = 32'b10011101101000000000000000000000;
    memory[49]   = 32'b01100010000000000000000000000000;
    memory[50]   = 32'b10011110001100000000000000000000;
    memory[51]   = 32'b00110000000000000000000000000000;
    memory[52]   = 32'b10011101101000000000000000000000;
    memory[53]   = 32'b10100000000000000000000000000000;
    memory[54]   = 32'b10100000000000000000000000000000;
    memory[55]   = 32'b11000110001010100000000000111100;
    memory[56]   = 32'b01011000000000000000000000000000;
    memory[57]   = 32'b01000000000000000000000000000000;
    memory[58]   = 32'b10000011000000000000000000000000;
    memory[59]   = 32'b11000000000000000000000000101010;
    memory[60]   = 32'b01011000000000000000000000000000;
    memory[61]   = 32'b01000000000000000000000000000000;
    memory[62]   = 32'b01110101000000000000000000000000;
    memory[63]   = 32'b01100010100000000000000000000000;
    memory[64]   = 32'b00111000000000000000000000000011;
    memory[65]   = 32'b01100100100000000000000000000000;
    memory[66]   = 32'b00111000000000000000000000000100;
    memory[67]   = 32'b01100101000000000000000000000000;
    memory[68]   = 32'b00100100000000000000000000000000;
    memory[69]   = 32'b11000000000000000000000001000110;
    memory[70]   = 32'b01010000000000000000000000000000;
    memory[71]   = 32'b00110000000000000000000000000000;
    memory[72]   = 32'b01011000000000000000000000000000;
    memory[73]   = 32'b01000000000000000000000000000000;
    memory[74]   = 32'b10000111000000000000000000000000;
    memory[75]   = 32'b11000100101010100000000001010110;
    memory[76]   = 32'b10000101000000000000000000000000;
    memory[77]   = 32'b11000100101010100000000001010110;
    memory[78]   = 32'b11000111001100100000000001010000;
    memory[79]   = 32'b11000000000000000000000001000101;
    memory[80]   = 32'b10011100101100000000000000000000;
    memory[81]   = 32'b00100100000000000000000000000000;
    memory[82]   = 32'b11110100100000000000000000000001;
    memory[83]   = 32'b11000100101010100000000001010110;
    memory[84]   = 32'b10000001000000000000000000000000;
    memory[85]   = 32'b11000000000000000000000001000110;
    memory[86]   = 32'b00011000000000000000000000000000;

	end
	
	always @(posedge clock) begin
	if (im_r==1)
		current_instruction <= memory[addr];
	else 
		current_instruction <= current_instruction;
	end
		
	assign instr_out = current_instruction;
endmodule	